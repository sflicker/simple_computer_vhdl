library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package Utils is
    function to_hex_string(byte : std_logic_vector(7 downto 0)) return string;

    
end Utils;